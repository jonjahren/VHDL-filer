library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity ghost_ram_lut is
   generic(
      ADDR_WIDTH : integer := 10;
      DATA_WIDTH : integer := 2
   );
   port(
      clk    : in  std_logic;
      we     : in  std_logic;
      addr_w : in  std_logic_vector(ADDR_WIDTH - 1 downto 0);
      addr_r : in  std_logic_vector(ADDR_WIDTH - 1 downto 0);
      din    : in  std_logic_vector(DATA_WIDTH - 1 downto 0);
      dout   : out std_logic_vector(DATA_WIDTH - 1 downto 0)
   );
end ghost_ram_lut;

architecture beh_arch of ghost_ram_lut is
   type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(DATA_WIDTH - 1 downto 0);
   -- sprite LUT
   constant INIT_GHOST_LUT : ram_type :=       
   (
      -- ghost sprite #0 
      "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
      "00", "00", "00", "00", "00", "00", "10", "10", "10", "10", "00", "00", "00", "00", "00", "00",
      "00", "00", "00", "00", "10", "10", "10", "10", "10", "10", "10", "10", "00", "00", "00", "00",
      "00", "00", "00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00", "00", "00",
      "00", "00", "00", "10", "10", "11", "11", "10", "10", "10", "10", "11", "11", "00", "00", "00",
      "00", "00", "10", "10", "11", "11", "11", "11", "10", "10", "11", "11", "11", "11", "00", "00",
      "00", "10", "10", "10", "11", "11", "01", "01", "10", "10", "11", "11", "01", "01", "00", "00",
      "00", "10", "10", "10", "11", "11", "01", "01", "10", "10", "11", "11", "01", "01", "10", "00",
      "00", "10", "10", "10", "10", "11", "11", "10", "10", "10", "10", "11", "11", "10", "10", "00",
      "00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00",
      "00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00",
      "00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00",
      "00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00",
      "00", "10", "10", "00", "10", "10", "10", "00", "00", "10", "10", "10", "00", "10", "10", "00",
      "00", "10", "00", "00", "00", "10", "10", "00", "00", "10", "10", "00", "00", "00", "10", "00",
      "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",

      -- ghost sprite #1 
      "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
      "00", "00", "00", "00", "00", "00", "10", "10", "10", "10", "00", "00", "00", "00", "00", "00",
      "00", "00", "00", "00", "10", "10", "10", "10", "10", "10", "10", "10", "00", "00", "00", "00",
      "00", "00", "00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00", "00", "00",
      "00", "00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00", "00",
      "00", "00", "10", "10", "11", "11", "10", "10", "10", "10", "11", "11", "10", "10", "00", "00",
      "00", "00", "10", "11", "11", "11", "11", "10", "10", "11", "11", "11", "11", "10", "00", "00",
      "00", "10", "10", "11", "11", "11", "11", "10", "10", "11", "11", "11", "11", "10", "10", "00",
      "00", "10", "10", "11", "01", "01", "11", "10", "10", "11", "01", "01", "11", "10", "10", "00",
      "00", "10", "10", "10", "01", "01", "10", "10", "10", "10", "01", "01", "10", "10", "10", "00",
      "00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00",
      "00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00",
      "00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00",
      "00", "10", "10", "10", "10", "00", "10", "10", "10", "10", "00", "10", "10", "10", "10", "00",
      "00", "00", "10", "10", "00", "00", "00", "10", "10", "00", "00", "00", "10", "10", "00", "00",
      "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",

      -- ghost sprite #2 
      "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
      "00", "00", "00", "00", "00", "00", "10", "10", "10", "10", "00", "00", "00", "00", "00", "00",
      "00", "00", "00", "00", "10", "10", "10", "10", "10", "10", "10", "10", "00", "00", "00", "00",
      "00", "00", "00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00", "00", "00",
      "00", "00", "10", "11", "11", "10", "10", "10", "10", "11", "11", "10", "10", "10", "00", "00",
      "00", "00", "11", "11", "11", "11", "10", "10", "11", "11", "11", "11", "10", "10", "00", "00",
      "00", "00", "01", "01", "11", "11", "10", "10", "01", "01", "11", "11", "10", "10", "00", "00",
      "00", "10", "01", "01", "11", "11", "10", "10", "01", "01", "11", "11", "10", "10", "10", "00",
      "00", "10", "10", "11", "11", "10", "10", "10", "10", "11", "11", "10", "10", "10", "10", "00",
      "00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00",
      "00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00",
      "00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00",
      "00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00",
      "00", "10", "10", "00", "10", "10", "10", "00", "00", "10", "10", "10", "00", "10", "10", "00",
      "00", "10", "00", "00", "00", "10", "10", "00", "00", "10", "10", "00", "00", "00", "10", "00",
      "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",

      -- ghost sprite #3 
      "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
      "00", "00", "00", "00", "00", "00", "10", "10", "10", "10", "00", "00", "00", "00", "00", "00",
      "00", "00", "00", "00", "01", "01", "10", "10", "10", "10", "01", "01", "00", "00", "00", "00",
      "00", "00", "00", "11", "01", "01", "11", "10", "10", "11", "01", "01", "11", "00", "00", "00",
      "00", "00", "10", "11", "11", "11", "11", "10", "10", "11", "11", "11", "11", "10", "00", "00",
      "00", "00", "10", "11", "11", "11", "11", "10", "10", "11", "11", "11", "11", "10", "00", "00",
      "00", "00", "10", "10", "11", "11", "10", "10", "10", "10", "11", "11", "10", "10", "00", "00",
      "00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00",
      "00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00",
      "00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00",
      "00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00",
      "00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00",
      "00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00",
      "00", "10", "10", "10", "10", "00", "10", "10", "10", "10", "00", "10", "10", "10", "10", "00",
      "00", "00", "10", "10", "00", "00", "00", "10", "10", "00", "00", "00", "10", "10", "00", "00",
      "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00"
   );
   signal ram : ram_type := INIT_GHOST_LUT;
begin
   process(clk)
   begin
      if (clk'event and clk = '1') then
         if (we = '1') then
            ram(to_integer(unsigned(addr_w))) <= din;
         end if;
         dout <= ram(to_integer(unsigned(addr_r)));
      end if;
   end process;
end beh_arch;
